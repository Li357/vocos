`timescale 1ns / 1ps
`default_nettype none

module mixer(
  input logic signed [31:0] carrier_channels  [N_FILTERS-1:0],
  input logic signed [31:0] envelope_channels [N_FILTERS-1:0],
);

  

endmodule

`default_nettype wire